----------------------------------------------------------------------------------
-- Company:    JHU EP
-- Engineer:   Ryan Newport
-- 
-- Create Date:   10/29/2018 
-- Module Name:   pwm
-- Project Name:  Lab06
--
-- Description:  pulse width modulation entity for mono-audio output signal
-----------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.all;

entity pwm is 
  Port()

