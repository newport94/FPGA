library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.all;


entity debounce is 
  Port(
    i_clk : in std_logic;
    i_rst : in std_logic);
end entity debounce;
  
architecture rtl of debounce is 

signal q_cntr

begin
  


end architecture rtl;
    